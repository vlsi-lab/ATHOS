module cbd (
    input athos_pkg::in_t cbd_i,
    input athos_pkg::funct7_t cycle_i, 
    output athos_pkg::out_t cbd_o
);

    logic [3:0] j;
    logic [31:0] d, a, b;
    logic [31:0] res;

    assign j = cbd_i.rs1_0[3:0];
    assign d = cbd_i.rs2_0;

    always_comb begin
        case(cycle_i.funct7_athos)
            athos_pkg::CBD3_1_MODE: begin
                a = d & 32'b00000000000000000000000000000111; //0x7
                b = {3'b000, d[31:3]} & 32'b00000000000000000000000000000111; //0x7
                res = a - b;
            end

            athos_pkg::CBD3_2_MODE: begin
                a = {6'b000000, d[31:6]} & 32'b00000000000000000000000000000111; //0x7
                b = {9'b000000000, d[31:9]} & 32'b00000000000000000000000000000111; //0x7
                res = a - b;
            end

            athos_pkg::CBD3_3_MODE: begin
                a = {12'b000000000000, d[31:12]} & 32'b00000000000000000000000000000111; //0x7
                b = {15'b000000000000000, d[31:15]} & 32'b00000000000000000000000000000111; //0x7
                res = a - b;
            end

            athos_pkg::CBD3_4_MODE: begin
                a = {18'b000000000000000000, d[31:18]} & 32'b00000000000000000000000000000111; //0x7
                b = {21'b000000000000000000000, d[31:21]} & 32'b00000000000000000000000000000111; //0x7
                res = a - b;
            end

            athos_pkg::CBD2_1_MODE: begin
                a = d & 32'b00000000000000000000000000000011; 
                b = {2'b00, d[31:2]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_2_MODE: begin
                a = {4'b0000 & d[31:4]} & 32'b00000000000000000000000000000011; 
                b = {6'b000000 & d[31:6]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_3_MODE: begin
                a = {8'b00000000 & d[31:8]} & 32'b00000000000000000000000000000011; 
                b = {10'b0000000000 & d[31:10]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_4_MODE: begin
                a = {12'b000000000000 & d[31:12]} & 32'b00000000000000000000000000000011; 
                b = {14'b00000000000000 & d[31:14]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_5_MODE: begin
                a = {16'b0000000000000000 & d[31:16]} & 32'b00000000000000000000000000000011; 
                b = {18'b000000000000000000 & d[31:18]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_6_MODE: begin
                a = {20'b00000000000000000000 & d[31:20]} & 32'b00000000000000000000000000000011; 
                b = {22'b0000000000000000000000 & d[31:22]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_7_MODE: begin
                a = {24'b000000000000000000000000 & d[31:24]} & 32'b00000000000000000000000000000011; 
                b = {26'b00000000000000000000000000 & d[31:26]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            athos_pkg::CBD2_8_MODE: begin
                a = {28'b0000000000000000000000000000 & d[31:28]} & 32'b00000000000000000000000000000011; 
                b = {30'b000000000000000000000000000000 & d[31:30]} & 32'b00000000000000000000000000000011; 
                res = a - b;
            end

            default: res = 'b0;  // Handle the default case if needed
        endcase
    end


    assign cbd_o.rd1 = '0;
    assign cbd_o.rd2 = res;

    
endmodule